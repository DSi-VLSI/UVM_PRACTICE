
class reg_transaction;
    
    base_pkg::ctrl_reg_t ctrl_reg;
    base_pkg::cfg_reg_t cfg_reg;
    base_pkg::clk_div_reg_t clk_div_reg;
    base_pkg::tx_fifo_stat_reg_t tx_fifo_stat_reg;
    base_pkg::rx_fifo_stat_reg_t rx_fifo_stat_reg;
    base_pkg::tx_fifo_data_reg_t tx_fifo_data_reg;
    base_pkg::rx_fifo_data_reg_t rx_fifo_data_reg;
    base_pkg::rx_fifo_peek_reg_t rx_fifo_peek_reg;

endclass