
package seq_pkg;

    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "define.svh"
    `include "seq_item.sv"
    `include "apb_base_seq.sv"
    `include "apb_write_seq.sv"
    `include "apb_read_seq.sv"
    `include "apb_reset_seq.sv"
    
endpackage