`include "axi/typedef.svh"

package base_pkg;

  `AXI_TYPEDEF_ALL(base, logic [31:0], logic [3:0], logic [63:0], logic [7:0], logic [7:0])

endpackage
