

interface uart_interface(input bit pclk);

    logic tx_o;
    logic rx_i;
    logic irq_o;
    
endinterface