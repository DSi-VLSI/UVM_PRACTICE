

interface uart_interface(input pclk);

    logic tx_o;
    logic rx_i;
    logic irq_o;
    
endinterface