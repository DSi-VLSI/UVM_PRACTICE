interface reset_intf
(
    input logic clk
);
    logic rst_n;
endinterface: reset_intf
