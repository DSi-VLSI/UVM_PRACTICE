

interface uart_interface();

    logic tx_o;
    logic rx_i;
    logic irq_o;
    
endinterface