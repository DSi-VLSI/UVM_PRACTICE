package environment_pkg;

    `include "uvm_macros.svh"
    import uvm_pkg::*;
    import seq_pkg::*;
    import apb_agent_pkg::*;
    import uart_agent_pkg::*;
    

    `include "uart_scoreboard.sv"
    `include "uart_environment.sv"
    
endpackage