`include "simple_test.sv"
`include "v_simple_test.sv"
