
package apb_agent_pkg;

    
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    import seq_pkg::*;

    `include "apb_sequencer.sv"
    `include "apb_driver.sv"
    `include "apb_monitor.sv"
    `include "apb_agent.sv"
    
    
endpackage