interface uart_intf(
    input  logic clk
);
    logic tx;
    logic rx;
    logic irq;
endinterface